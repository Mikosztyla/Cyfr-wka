library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fpga is
	port (
		clk : in std_logic;
		spd_input : in std_logic;
		rvs_input : in std_logic;
		left_out : out std_logic_vector(7 downto 0);
		right_out : out std_logic_vector(7 downto 0)
	);
end fpga;


architecture snake of fpga is
	signal state : unsigned(2 downto 0) := b"000";
	
	signal reverse_state: std_logic := '0';
	signal speed_state: std_logic := '0';

	constant fast_delay : integer := 10_000_000;
	constant slow_delay : integer := 3 * fast_delay;
	signal delay : integer := slow_delay;
	signal clock_counter : integer range 0 to 40_000_000;
	
	signal spd_input_history : std_logic_vector(7 downto 0) := (others => '0');
    signal rvs_input_history : std_logic_vector(7 downto 0) := (others => '0');

	begin
	
	SPEED : process(spd_input)
	begin
		spd_input_history <= spd_input_history(6 downto 0) & spd_input;
		if spd_input_history = "11111111" then
			if speed_state = '1' then
				speed_state <= '0';
				delay <= slow_delay;
			else
				speed_state <= '1';
				delay <= fast_delay;
			end if;
		end if;
	end process SPEED;
	
	DIRECTION : process(rvs_input)
	begin
		rvs_input_history <= rvs_input_history(6 downto 0) & rvs_input;
		if rvs_input_history = "11111111" then
			if reverse_state = '0' then
				reverse_state <= '1';
			else
				reverse_state <= '0';
			end if;
		end if;
	end process DIRECTION;

	
	MOVE: process(clk)
	begin
		if clk = '1' then
			clock_counter <= clock_counter + 1;
			
			if clock_counter >= delay then
				if reverse_state = '0' then
					state <= state + 1;
				else
					state <= state -1;
				end if;
				
				clock_counter <= 0;
			end if;
		end if;
	end process MOVE;
	
	
	DISPLAY : process(state)
	begin
		case state is
		when "000" => 
			left_out <= b"11110111";
			right_out <= b"11110111";
		when "001" => 
			left_out <= b"11111111";
			right_out <= b"11110011";
		when "010" => 
			left_out <= b"11111111";
			right_out <= b"11111001";
		when "011" => 
			left_out <= b"11111111";
			right_out <= b"10111101";
		when "100" => 
			left_out <= b"10111111";
			right_out <= b"10111111";
		when "101" => 
			left_out <= b"10011111";
			right_out <= b"11111111";
		when "110" => 
			left_out <= b"11001111";
			right_out <= b"11111111";
		when "111" => 
			left_out <= b"11100111";
			right_out <= b"11111111";
		when others =>
			left_out <= b"11111111";
			right_out <= b"11111111";
		end case;
		
	end process DISPLAY;
		
end snake;	
	